/*
 * id: 5
 * logic_id: 0
 * name: 输出0
 * level: 1
 * tags: 
 * points: 1
 */

module Zero(
    output out
);
    // 在这里输入你的代码 请不要修改模块和信号名称
    assign out = 0;
endmodule
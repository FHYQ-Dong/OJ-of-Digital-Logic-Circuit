/*
 * id: 6
 * logic_id: 1
 * name: 输出1
 * level: 1
 * tags: 
 * points: 1
 */

module One(
    output out
);
    // 在这里输入你的代码 请不要修改模块和信号名称
    assign out = 1;
endmodule